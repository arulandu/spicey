.title Voltage Divider
R1 in out 9k
R2 out in 1.5E-2
R3 in out 100Ohm
.end