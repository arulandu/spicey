.title Empty
.end